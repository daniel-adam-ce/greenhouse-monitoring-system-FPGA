// nios_system.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module nios_system (
		output wire        bme_csn_export,     //     bme_csn.export
		input  wire        bme_irq_export,     //     bme_irq.export
		input  wire        bme_miso_export,    //    bme_miso.export
		output wire        bme_mosi_export,    //    bme_mosi.export
		output wire        bme_sck_export,     //     bme_sck.export
		input  wire        clk_clk,            //         clk.clk
		input  wire [3:0]  keys_export,        //        keys.export
		output wire [7:0]  leds_g_export,      //      leds_g.export
		output wire [31:0] leds_r_export,      //      leds_r.export
		output wire        nrf_ce_export,      //      nrf_ce.export
		output wire        nrf_csn_export,     //     nrf_csn.export
		input  wire        nrf_irq_export,     //     nrf_irq.export
		input  wire        nrf_miso_export,    //    nrf_miso.export
		output wire        nrf_mosi_export,    //    nrf_mosi.export
		output wire        nrf_sck_export,     //     nrf_sck.export
		input  wire        reset_reset,        //       reset.reset
		output wire [11:0] sdram_addr,         //       sdram.addr
		output wire [1:0]  sdram_ba,           //            .ba
		output wire        sdram_cas_n,        //            .cas_n
		output wire        sdram_cke,          //            .cke
		output wire        sdram_cs_n,         //            .cs_n
		inout  wire [31:0] sdram_dq,           //            .dq
		output wire [3:0]  sdram_dqm,          //            .dqm
		output wire        sdram_ras_n,        //            .ras_n
		output wire        sdram_we_n,         //            .we_n
		output wire        sdram_clk_clk,      //   sdram_clk.clk
		output wire [31:0] seven_seg_0_export, // seven_seg_0.export
		output wire [31:0] seven_seg_1_export, // seven_seg_1.export
		input  wire [31:0] switches_export     //    switches.export
	);

	wire         sys_sdram_pll_0_sys_clk_clk;                                 // sys_sdram_pll_0:sys_clk_clk -> [bme_csn:clk, bme_irq:clk, bme_miso:clk, bme_mosi:clk, bme_sck:clk, irq_mapper:clk, jtag_uart_0:clk, keys:clk, leds_g:clk, leds_r:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, new_sdram_controller_0:clk, nios2_gen2_0:clk, nrf_ce:clk, nrf_csn:clk, nrf_irq:clk, nrf_miso:clk, nrf_mosi:clk, nrf_sck:clk, onchip_memory2_0:clk, rst_controller:clk, seven_seg_0:clk, seven_seg_1:clk, switches:clk, sysid_qsys_0:clock, timer_0:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                      // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                       // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_leds_r_s1_chipselect;                      // mm_interconnect_0:leds_r_s1_chipselect -> leds_r:chipselect
	wire  [31:0] mm_interconnect_0_leds_r_s1_readdata;                        // leds_r:readdata -> mm_interconnect_0:leds_r_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_r_s1_address;                         // mm_interconnect_0:leds_r_s1_address -> leds_r:address
	wire         mm_interconnect_0_leds_r_s1_write;                           // mm_interconnect_0:leds_r_s1_write -> leds_r:write_n
	wire  [31:0] mm_interconnect_0_leds_r_s1_writedata;                       // mm_interconnect_0:leds_r_s1_writedata -> leds_r:writedata
	wire         mm_interconnect_0_seven_seg_0_s1_chipselect;                 // mm_interconnect_0:seven_seg_0_s1_chipselect -> seven_seg_0:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_0_s1_readdata;                   // seven_seg_0:readdata -> mm_interconnect_0:seven_seg_0_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_0_s1_address;                    // mm_interconnect_0:seven_seg_0_s1_address -> seven_seg_0:address
	wire         mm_interconnect_0_seven_seg_0_s1_write;                      // mm_interconnect_0:seven_seg_0_s1_write -> seven_seg_0:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_0_s1_writedata;                  // mm_interconnect_0:seven_seg_0_s1_writedata -> seven_seg_0:writedata
	wire         mm_interconnect_0_seven_seg_1_s1_chipselect;                 // mm_interconnect_0:seven_seg_1_s1_chipselect -> seven_seg_1:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_1_s1_readdata;                   // seven_seg_1:readdata -> mm_interconnect_0:seven_seg_1_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_1_s1_address;                    // mm_interconnect_0:seven_seg_1_s1_address -> seven_seg_1:address
	wire         mm_interconnect_0_seven_seg_1_s1_write;                      // mm_interconnect_0:seven_seg_1_s1_write -> seven_seg_1:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_1_s1_writedata;                  // mm_interconnect_0:seven_seg_1_s1_writedata -> seven_seg_1:writedata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_chipselect;      // mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire  [31:0] mm_interconnect_0_new_sdram_controller_0_s1_readdata;        // new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_waitrequest;     // new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	wire  [21:0] mm_interconnect_0_new_sdram_controller_0_s1_address;         // mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire         mm_interconnect_0_new_sdram_controller_0_s1_read;            // mm_interconnect_0:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire   [3:0] mm_interconnect_0_new_sdram_controller_0_s1_byteenable;      // mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire         mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid;   // new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_0_new_sdram_controller_0_s1_write;           // mm_interconnect_0:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire  [31:0] mm_interconnect_0_new_sdram_controller_0_s1_writedata;       // mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire         mm_interconnect_0_keys_s1_chipselect;                        // mm_interconnect_0:keys_s1_chipselect -> keys:chipselect
	wire  [31:0] mm_interconnect_0_keys_s1_readdata;                          // keys:readdata -> mm_interconnect_0:keys_s1_readdata
	wire   [1:0] mm_interconnect_0_keys_s1_address;                           // mm_interconnect_0:keys_s1_address -> keys:address
	wire         mm_interconnect_0_keys_s1_write;                             // mm_interconnect_0:keys_s1_write -> keys:write_n
	wire  [31:0] mm_interconnect_0_keys_s1_writedata;                         // mm_interconnect_0:keys_s1_writedata -> keys:writedata
	wire         mm_interconnect_0_leds_g_s1_chipselect;                      // mm_interconnect_0:leds_g_s1_chipselect -> leds_g:chipselect
	wire  [31:0] mm_interconnect_0_leds_g_s1_readdata;                        // leds_g:readdata -> mm_interconnect_0:leds_g_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_g_s1_address;                         // mm_interconnect_0:leds_g_s1_address -> leds_g:address
	wire         mm_interconnect_0_leds_g_s1_write;                           // mm_interconnect_0:leds_g_s1_write -> leds_g:write_n
	wire  [31:0] mm_interconnect_0_leds_g_s1_writedata;                       // mm_interconnect_0:leds_g_s1_writedata -> leds_g:writedata
	wire         mm_interconnect_0_bme_csn_s1_chipselect;                     // mm_interconnect_0:bme_csn_s1_chipselect -> bme_csn:chipselect
	wire  [31:0] mm_interconnect_0_bme_csn_s1_readdata;                       // bme_csn:readdata -> mm_interconnect_0:bme_csn_s1_readdata
	wire   [1:0] mm_interconnect_0_bme_csn_s1_address;                        // mm_interconnect_0:bme_csn_s1_address -> bme_csn:address
	wire         mm_interconnect_0_bme_csn_s1_write;                          // mm_interconnect_0:bme_csn_s1_write -> bme_csn:write_n
	wire  [31:0] mm_interconnect_0_bme_csn_s1_writedata;                      // mm_interconnect_0:bme_csn_s1_writedata -> bme_csn:writedata
	wire         mm_interconnect_0_bme_sck_s1_chipselect;                     // mm_interconnect_0:bme_sck_s1_chipselect -> bme_sck:chipselect
	wire  [31:0] mm_interconnect_0_bme_sck_s1_readdata;                       // bme_sck:readdata -> mm_interconnect_0:bme_sck_s1_readdata
	wire   [1:0] mm_interconnect_0_bme_sck_s1_address;                        // mm_interconnect_0:bme_sck_s1_address -> bme_sck:address
	wire         mm_interconnect_0_bme_sck_s1_write;                          // mm_interconnect_0:bme_sck_s1_write -> bme_sck:write_n
	wire  [31:0] mm_interconnect_0_bme_sck_s1_writedata;                      // mm_interconnect_0:bme_sck_s1_writedata -> bme_sck:writedata
	wire         mm_interconnect_0_bme_mosi_s1_chipselect;                    // mm_interconnect_0:bme_mosi_s1_chipselect -> bme_mosi:chipselect
	wire  [31:0] mm_interconnect_0_bme_mosi_s1_readdata;                      // bme_mosi:readdata -> mm_interconnect_0:bme_mosi_s1_readdata
	wire   [1:0] mm_interconnect_0_bme_mosi_s1_address;                       // mm_interconnect_0:bme_mosi_s1_address -> bme_mosi:address
	wire         mm_interconnect_0_bme_mosi_s1_write;                         // mm_interconnect_0:bme_mosi_s1_write -> bme_mosi:write_n
	wire  [31:0] mm_interconnect_0_bme_mosi_s1_writedata;                     // mm_interconnect_0:bme_mosi_s1_writedata -> bme_mosi:writedata
	wire  [31:0] mm_interconnect_0_bme_miso_s1_readdata;                      // bme_miso:readdata -> mm_interconnect_0:bme_miso_s1_readdata
	wire   [1:0] mm_interconnect_0_bme_miso_s1_address;                       // mm_interconnect_0:bme_miso_s1_address -> bme_miso:address
	wire         mm_interconnect_0_bme_irq_s1_chipselect;                     // mm_interconnect_0:bme_irq_s1_chipselect -> bme_irq:chipselect
	wire  [31:0] mm_interconnect_0_bme_irq_s1_readdata;                       // bme_irq:readdata -> mm_interconnect_0:bme_irq_s1_readdata
	wire   [1:0] mm_interconnect_0_bme_irq_s1_address;                        // mm_interconnect_0:bme_irq_s1_address -> bme_irq:address
	wire         mm_interconnect_0_bme_irq_s1_write;                          // mm_interconnect_0:bme_irq_s1_write -> bme_irq:write_n
	wire  [31:0] mm_interconnect_0_bme_irq_s1_writedata;                      // mm_interconnect_0:bme_irq_s1_writedata -> bme_irq:writedata
	wire         mm_interconnect_0_nrf_csn_s1_chipselect;                     // mm_interconnect_0:nrf_csn_s1_chipselect -> nrf_csn:chipselect
	wire  [31:0] mm_interconnect_0_nrf_csn_s1_readdata;                       // nrf_csn:readdata -> mm_interconnect_0:nrf_csn_s1_readdata
	wire   [1:0] mm_interconnect_0_nrf_csn_s1_address;                        // mm_interconnect_0:nrf_csn_s1_address -> nrf_csn:address
	wire         mm_interconnect_0_nrf_csn_s1_write;                          // mm_interconnect_0:nrf_csn_s1_write -> nrf_csn:write_n
	wire  [31:0] mm_interconnect_0_nrf_csn_s1_writedata;                      // mm_interconnect_0:nrf_csn_s1_writedata -> nrf_csn:writedata
	wire         mm_interconnect_0_nrf_sck_s1_chipselect;                     // mm_interconnect_0:nrf_sck_s1_chipselect -> nrf_sck:chipselect
	wire  [31:0] mm_interconnect_0_nrf_sck_s1_readdata;                       // nrf_sck:readdata -> mm_interconnect_0:nrf_sck_s1_readdata
	wire   [1:0] mm_interconnect_0_nrf_sck_s1_address;                        // mm_interconnect_0:nrf_sck_s1_address -> nrf_sck:address
	wire         mm_interconnect_0_nrf_sck_s1_write;                          // mm_interconnect_0:nrf_sck_s1_write -> nrf_sck:write_n
	wire  [31:0] mm_interconnect_0_nrf_sck_s1_writedata;                      // mm_interconnect_0:nrf_sck_s1_writedata -> nrf_sck:writedata
	wire         mm_interconnect_0_nrf_mosi_s1_chipselect;                    // mm_interconnect_0:nrf_mosi_s1_chipselect -> nrf_mosi:chipselect
	wire  [31:0] mm_interconnect_0_nrf_mosi_s1_readdata;                      // nrf_mosi:readdata -> mm_interconnect_0:nrf_mosi_s1_readdata
	wire   [1:0] mm_interconnect_0_nrf_mosi_s1_address;                       // mm_interconnect_0:nrf_mosi_s1_address -> nrf_mosi:address
	wire         mm_interconnect_0_nrf_mosi_s1_write;                         // mm_interconnect_0:nrf_mosi_s1_write -> nrf_mosi:write_n
	wire  [31:0] mm_interconnect_0_nrf_mosi_s1_writedata;                     // mm_interconnect_0:nrf_mosi_s1_writedata -> nrf_mosi:writedata
	wire  [31:0] mm_interconnect_0_nrf_miso_s1_readdata;                      // nrf_miso:readdata -> mm_interconnect_0:nrf_miso_s1_readdata
	wire   [1:0] mm_interconnect_0_nrf_miso_s1_address;                       // mm_interconnect_0:nrf_miso_s1_address -> nrf_miso:address
	wire         mm_interconnect_0_nrf_ce_s1_chipselect;                      // mm_interconnect_0:nrf_ce_s1_chipselect -> nrf_ce:chipselect
	wire  [31:0] mm_interconnect_0_nrf_ce_s1_readdata;                        // nrf_ce:readdata -> mm_interconnect_0:nrf_ce_s1_readdata
	wire   [1:0] mm_interconnect_0_nrf_ce_s1_address;                         // mm_interconnect_0:nrf_ce_s1_address -> nrf_ce:address
	wire         mm_interconnect_0_nrf_ce_s1_write;                           // mm_interconnect_0:nrf_ce_s1_write -> nrf_ce:write_n
	wire  [31:0] mm_interconnect_0_nrf_ce_s1_writedata;                       // mm_interconnect_0:nrf_ce_s1_writedata -> nrf_ce:writedata
	wire         mm_interconnect_0_nrf_irq_s1_chipselect;                     // mm_interconnect_0:nrf_irq_s1_chipselect -> nrf_irq:chipselect
	wire  [31:0] mm_interconnect_0_nrf_irq_s1_readdata;                       // nrf_irq:readdata -> mm_interconnect_0:nrf_irq_s1_readdata
	wire   [1:0] mm_interconnect_0_nrf_irq_s1_address;                        // mm_interconnect_0:nrf_irq_s1_address -> nrf_irq:address
	wire         mm_interconnect_0_nrf_irq_s1_write;                          // mm_interconnect_0:nrf_irq_s1_write -> nrf_irq:write_n
	wire  [31:0] mm_interconnect_0_nrf_irq_s1_writedata;                      // mm_interconnect_0:nrf_irq_s1_writedata -> nrf_irq:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // keys:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // bme_irq:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                    // nrf_irq:irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [bme_csn:reset_n, bme_irq:reset_n, bme_miso:reset_n, bme_mosi:reset_n, bme_sck:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, keys:reset_n, leds_g:reset_n, leds_r:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n, nios2_gen2_0:reset_n, nrf_ce:reset_n, nrf_csn:reset_n, nrf_irq:reset_n, nrf_miso:reset_n, nrf_mosi:reset_n, nrf_sck:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, seven_seg_0:reset_n, seven_seg_1:reset_n, switches:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> rst_controller:reset_in0

	nios_system_bme_csn bme_csn (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_bme_csn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bme_csn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bme_csn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bme_csn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bme_csn_s1_readdata),   //                    .readdata
		.out_port   (bme_csn_export)                           // external_connection.export
	);

	nios_system_bme_irq bme_irq (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_bme_irq_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bme_irq_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bme_irq_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bme_irq_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bme_irq_s1_readdata),   //                    .readdata
		.in_port    (bme_irq_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                 //                 irq.irq
	);

	nios_system_bme_miso bme_miso (
		.clk      (sys_sdram_pll_0_sys_clk_clk),            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_bme_miso_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_bme_miso_s1_readdata), //                    .readdata
		.in_port  (bme_miso_export)                         // external_connection.export
	);

	nios_system_bme_csn bme_mosi (
		.clk        (sys_sdram_pll_0_sys_clk_clk),              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bme_mosi_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bme_mosi_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bme_mosi_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bme_mosi_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bme_mosi_s1_readdata),   //                    .readdata
		.out_port   (bme_mosi_export)                           // external_connection.export
	);

	nios_system_bme_csn bme_sck (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_bme_sck_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bme_sck_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bme_sck_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bme_sck_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bme_sck_s1_readdata),   //                    .readdata
		.out_port   (bme_sck_export)                           // external_connection.export
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                                 //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_keys keys (
		.clk        (sys_sdram_pll_0_sys_clk_clk),          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_keys_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keys_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keys_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keys_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keys_s1_readdata),   //                    .readdata
		.in_port    (keys_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)              //                 irq.irq
	);

	nios_system_leds_g leds_g (
		.clk        (sys_sdram_pll_0_sys_clk_clk),            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_leds_g_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_g_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_g_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_g_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_g_s1_readdata),   //                    .readdata
		.out_port   (leds_g_export)                           // external_connection.export
	);

	nios_system_leds_r leds_r (
		.clk        (sys_sdram_pll_0_sys_clk_clk),            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_leds_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_r_s1_readdata),   //                    .readdata
		.out_port   (leds_r_export)                           // external_connection.export
	);

	nios_system_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                           // reset.reset_n
		.az_addr        (mm_interconnect_0_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                                //  wire.export
		.zs_ba          (sdram_ba),                                                  //      .export
		.zs_cas_n       (sdram_cas_n),                                               //      .export
		.zs_cke         (sdram_cke),                                                 //      .export
		.zs_cs_n        (sdram_cs_n),                                                //      .export
		.zs_dq          (sdram_dq),                                                  //      .export
		.zs_dqm         (sdram_dqm),                                                 //      .export
		.zs_ras_n       (sdram_ras_n),                                               //      .export
		.zs_we_n        (sdram_we_n)                                                 //      .export
	);

	nios_system_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (sys_sdram_pll_0_sys_clk_clk),                                //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_system_bme_csn nrf_ce (
		.clk        (sys_sdram_pll_0_sys_clk_clk),            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_nrf_ce_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nrf_ce_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nrf_ce_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nrf_ce_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nrf_ce_s1_readdata),   //                    .readdata
		.out_port   (nrf_ce_export)                           // external_connection.export
	);

	nios_system_bme_csn nrf_csn (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_nrf_csn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nrf_csn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nrf_csn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nrf_csn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nrf_csn_s1_readdata),   //                    .readdata
		.out_port   (nrf_csn_export)                           // external_connection.export
	);

	nios_system_bme_irq nrf_irq (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_nrf_irq_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nrf_irq_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nrf_irq_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nrf_irq_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nrf_irq_s1_readdata),   //                    .readdata
		.in_port    (nrf_irq_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                 //                 irq.irq
	);

	nios_system_bme_miso nrf_miso (
		.clk      (sys_sdram_pll_0_sys_clk_clk),            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_nrf_miso_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_nrf_miso_s1_readdata), //                    .readdata
		.in_port  (nrf_miso_export)                         // external_connection.export
	);

	nios_system_bme_csn nrf_mosi (
		.clk        (sys_sdram_pll_0_sys_clk_clk),              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_nrf_mosi_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nrf_mosi_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nrf_mosi_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nrf_mosi_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nrf_mosi_s1_readdata),   //                    .readdata
		.out_port   (nrf_mosi_export)                           // external_connection.export
	);

	nios_system_bme_csn nrf_sck (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_nrf_sck_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nrf_sck_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nrf_sck_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nrf_sck_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nrf_sck_s1_readdata),   //                    .readdata
		.out_port   (nrf_sck_export)                           // external_connection.export
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                      //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	nios_system_leds_r seven_seg_0 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_0_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_0_export)                           // external_connection.export
	);

	nios_system_leds_r seven_seg_1 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_1_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_1_export)                           // external_connection.export
	);

	nios_system_switches switches (
		.clk      (sys_sdram_pll_0_sys_clk_clk),            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	nios_system_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (clk_clk),                     //      ref_clk.clk
		.ref_reset_reset    (reset_reset),                 //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_0_sys_clk_clk), //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),               //    sdram_clk.clk
		.reset_source_reset ()                             // reset_source.reset
	);

	nios_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (sys_sdram_pll_0_sys_clk_clk),                           //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_system_timer_0 timer_0 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),             //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.sys_sdram_pll_0_sys_clk_clk                    (sys_sdram_pll_0_sys_clk_clk),                                 //                  sys_sdram_pll_0_sys_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_readdatavalid         (nios2_gen2_0_data_master_readdatavalid),                      //                                         .readdatavalid
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.nios2_gen2_0_instruction_master_readdatavalid  (nios2_gen2_0_instruction_master_readdatavalid),               //                                         .readdatavalid
		.bme_csn_s1_address                             (mm_interconnect_0_bme_csn_s1_address),                        //                               bme_csn_s1.address
		.bme_csn_s1_write                               (mm_interconnect_0_bme_csn_s1_write),                          //                                         .write
		.bme_csn_s1_readdata                            (mm_interconnect_0_bme_csn_s1_readdata),                       //                                         .readdata
		.bme_csn_s1_writedata                           (mm_interconnect_0_bme_csn_s1_writedata),                      //                                         .writedata
		.bme_csn_s1_chipselect                          (mm_interconnect_0_bme_csn_s1_chipselect),                     //                                         .chipselect
		.bme_irq_s1_address                             (mm_interconnect_0_bme_irq_s1_address),                        //                               bme_irq_s1.address
		.bme_irq_s1_write                               (mm_interconnect_0_bme_irq_s1_write),                          //                                         .write
		.bme_irq_s1_readdata                            (mm_interconnect_0_bme_irq_s1_readdata),                       //                                         .readdata
		.bme_irq_s1_writedata                           (mm_interconnect_0_bme_irq_s1_writedata),                      //                                         .writedata
		.bme_irq_s1_chipselect                          (mm_interconnect_0_bme_irq_s1_chipselect),                     //                                         .chipselect
		.bme_miso_s1_address                            (mm_interconnect_0_bme_miso_s1_address),                       //                              bme_miso_s1.address
		.bme_miso_s1_readdata                           (mm_interconnect_0_bme_miso_s1_readdata),                      //                                         .readdata
		.bme_mosi_s1_address                            (mm_interconnect_0_bme_mosi_s1_address),                       //                              bme_mosi_s1.address
		.bme_mosi_s1_write                              (mm_interconnect_0_bme_mosi_s1_write),                         //                                         .write
		.bme_mosi_s1_readdata                           (mm_interconnect_0_bme_mosi_s1_readdata),                      //                                         .readdata
		.bme_mosi_s1_writedata                          (mm_interconnect_0_bme_mosi_s1_writedata),                     //                                         .writedata
		.bme_mosi_s1_chipselect                         (mm_interconnect_0_bme_mosi_s1_chipselect),                    //                                         .chipselect
		.bme_sck_s1_address                             (mm_interconnect_0_bme_sck_s1_address),                        //                               bme_sck_s1.address
		.bme_sck_s1_write                               (mm_interconnect_0_bme_sck_s1_write),                          //                                         .write
		.bme_sck_s1_readdata                            (mm_interconnect_0_bme_sck_s1_readdata),                       //                                         .readdata
		.bme_sck_s1_writedata                           (mm_interconnect_0_bme_sck_s1_writedata),                      //                                         .writedata
		.bme_sck_s1_chipselect                          (mm_interconnect_0_bme_sck_s1_chipselect),                     //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.keys_s1_address                                (mm_interconnect_0_keys_s1_address),                           //                                  keys_s1.address
		.keys_s1_write                                  (mm_interconnect_0_keys_s1_write),                             //                                         .write
		.keys_s1_readdata                               (mm_interconnect_0_keys_s1_readdata),                          //                                         .readdata
		.keys_s1_writedata                              (mm_interconnect_0_keys_s1_writedata),                         //                                         .writedata
		.keys_s1_chipselect                             (mm_interconnect_0_keys_s1_chipselect),                        //                                         .chipselect
		.leds_g_s1_address                              (mm_interconnect_0_leds_g_s1_address),                         //                                leds_g_s1.address
		.leds_g_s1_write                                (mm_interconnect_0_leds_g_s1_write),                           //                                         .write
		.leds_g_s1_readdata                             (mm_interconnect_0_leds_g_s1_readdata),                        //                                         .readdata
		.leds_g_s1_writedata                            (mm_interconnect_0_leds_g_s1_writedata),                       //                                         .writedata
		.leds_g_s1_chipselect                           (mm_interconnect_0_leds_g_s1_chipselect),                      //                                         .chipselect
		.leds_r_s1_address                              (mm_interconnect_0_leds_r_s1_address),                         //                                leds_r_s1.address
		.leds_r_s1_write                                (mm_interconnect_0_leds_r_s1_write),                           //                                         .write
		.leds_r_s1_readdata                             (mm_interconnect_0_leds_r_s1_readdata),                        //                                         .readdata
		.leds_r_s1_writedata                            (mm_interconnect_0_leds_r_s1_writedata),                       //                                         .writedata
		.leds_r_s1_chipselect                           (mm_interconnect_0_leds_r_s1_chipselect),                      //                                         .chipselect
		.new_sdram_controller_0_s1_address              (mm_interconnect_0_new_sdram_controller_0_s1_address),         //                new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write                (mm_interconnect_0_new_sdram_controller_0_s1_write),           //                                         .write
		.new_sdram_controller_0_s1_read                 (mm_interconnect_0_new_sdram_controller_0_s1_read),            //                                         .read
		.new_sdram_controller_0_s1_readdata             (mm_interconnect_0_new_sdram_controller_0_s1_readdata),        //                                         .readdata
		.new_sdram_controller_0_s1_writedata            (mm_interconnect_0_new_sdram_controller_0_s1_writedata),       //                                         .writedata
		.new_sdram_controller_0_s1_byteenable           (mm_interconnect_0_new_sdram_controller_0_s1_byteenable),      //                                         .byteenable
		.new_sdram_controller_0_s1_readdatavalid        (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid),   //                                         .readdatavalid
		.new_sdram_controller_0_s1_waitrequest          (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),     //                                         .waitrequest
		.new_sdram_controller_0_s1_chipselect           (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),      //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.nrf_ce_s1_address                              (mm_interconnect_0_nrf_ce_s1_address),                         //                                nrf_ce_s1.address
		.nrf_ce_s1_write                                (mm_interconnect_0_nrf_ce_s1_write),                           //                                         .write
		.nrf_ce_s1_readdata                             (mm_interconnect_0_nrf_ce_s1_readdata),                        //                                         .readdata
		.nrf_ce_s1_writedata                            (mm_interconnect_0_nrf_ce_s1_writedata),                       //                                         .writedata
		.nrf_ce_s1_chipselect                           (mm_interconnect_0_nrf_ce_s1_chipselect),                      //                                         .chipselect
		.nrf_csn_s1_address                             (mm_interconnect_0_nrf_csn_s1_address),                        //                               nrf_csn_s1.address
		.nrf_csn_s1_write                               (mm_interconnect_0_nrf_csn_s1_write),                          //                                         .write
		.nrf_csn_s1_readdata                            (mm_interconnect_0_nrf_csn_s1_readdata),                       //                                         .readdata
		.nrf_csn_s1_writedata                           (mm_interconnect_0_nrf_csn_s1_writedata),                      //                                         .writedata
		.nrf_csn_s1_chipselect                          (mm_interconnect_0_nrf_csn_s1_chipselect),                     //                                         .chipselect
		.nrf_irq_s1_address                             (mm_interconnect_0_nrf_irq_s1_address),                        //                               nrf_irq_s1.address
		.nrf_irq_s1_write                               (mm_interconnect_0_nrf_irq_s1_write),                          //                                         .write
		.nrf_irq_s1_readdata                            (mm_interconnect_0_nrf_irq_s1_readdata),                       //                                         .readdata
		.nrf_irq_s1_writedata                           (mm_interconnect_0_nrf_irq_s1_writedata),                      //                                         .writedata
		.nrf_irq_s1_chipselect                          (mm_interconnect_0_nrf_irq_s1_chipselect),                     //                                         .chipselect
		.nrf_miso_s1_address                            (mm_interconnect_0_nrf_miso_s1_address),                       //                              nrf_miso_s1.address
		.nrf_miso_s1_readdata                           (mm_interconnect_0_nrf_miso_s1_readdata),                      //                                         .readdata
		.nrf_mosi_s1_address                            (mm_interconnect_0_nrf_mosi_s1_address),                       //                              nrf_mosi_s1.address
		.nrf_mosi_s1_write                              (mm_interconnect_0_nrf_mosi_s1_write),                         //                                         .write
		.nrf_mosi_s1_readdata                           (mm_interconnect_0_nrf_mosi_s1_readdata),                      //                                         .readdata
		.nrf_mosi_s1_writedata                          (mm_interconnect_0_nrf_mosi_s1_writedata),                     //                                         .writedata
		.nrf_mosi_s1_chipselect                         (mm_interconnect_0_nrf_mosi_s1_chipselect),                    //                                         .chipselect
		.nrf_sck_s1_address                             (mm_interconnect_0_nrf_sck_s1_address),                        //                               nrf_sck_s1.address
		.nrf_sck_s1_write                               (mm_interconnect_0_nrf_sck_s1_write),                          //                                         .write
		.nrf_sck_s1_readdata                            (mm_interconnect_0_nrf_sck_s1_readdata),                       //                                         .readdata
		.nrf_sck_s1_writedata                           (mm_interconnect_0_nrf_sck_s1_writedata),                      //                                         .writedata
		.nrf_sck_s1_chipselect                          (mm_interconnect_0_nrf_sck_s1_chipselect),                     //                                         .chipselect
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.seven_seg_0_s1_address                         (mm_interconnect_0_seven_seg_0_s1_address),                    //                           seven_seg_0_s1.address
		.seven_seg_0_s1_write                           (mm_interconnect_0_seven_seg_0_s1_write),                      //                                         .write
		.seven_seg_0_s1_readdata                        (mm_interconnect_0_seven_seg_0_s1_readdata),                   //                                         .readdata
		.seven_seg_0_s1_writedata                       (mm_interconnect_0_seven_seg_0_s1_writedata),                  //                                         .writedata
		.seven_seg_0_s1_chipselect                      (mm_interconnect_0_seven_seg_0_s1_chipselect),                 //                                         .chipselect
		.seven_seg_1_s1_address                         (mm_interconnect_0_seven_seg_1_s1_address),                    //                           seven_seg_1_s1.address
		.seven_seg_1_s1_write                           (mm_interconnect_0_seven_seg_1_s1_write),                      //                                         .write
		.seven_seg_1_s1_readdata                        (mm_interconnect_0_seven_seg_1_s1_readdata),                   //                                         .readdata
		.seven_seg_1_s1_writedata                       (mm_interconnect_0_seven_seg_1_s1_writedata),                  //                                         .writedata
		.seven_seg_1_s1_chipselect                      (mm_interconnect_0_seven_seg_1_s1_chipselect),                 //                                         .chipselect
		.switches_s1_address                            (mm_interconnect_0_switches_s1_address),                       //                              switches_s1.address
		.switches_s1_readdata                           (mm_interconnect_0_switches_s1_readdata),                      //                                         .readdata
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                         .readdata
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                        //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                          //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                       //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                      //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect)                      //                                         .chipselect
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (sys_sdram_pll_0_sys_clk_clk),    //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
